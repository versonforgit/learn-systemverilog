module test(input clk_i,
            input rstn_i,
            input [1:0] cmd_i,
            output [1:0] slv0_prio,
            output [2:0] slv0_len,
            output [1:0] slv_o);
endmodule